`ifndef AXI_PKG_SVH_
`define AXI_PKG_SVH_

package axi_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "axi_define.svh"
`include "axi_trans.svh"
`include "axi_sequencer.svh"
`include "axi_slv_driver.svh"
`include "axi_monitor.svh"
`include "axi_agent.svh"

endpackage : axi_pkg
`endif
