`ifndef AHB_PKG_SVH_
`define AHB_PKG_SVH_

package ahb_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "ahb_type.svh"
`include "ahb_trans.svh"
`include "ahb_sequencer.svh"
`include "ahb_master_driver.svh"
`include "ahb_monitor.svh"
`include "ahb_agent.svh"
`include "ahb_adapter.svh"

endpackage : ahb_pkg
`endif
